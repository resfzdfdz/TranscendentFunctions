/*******************************************************************************
  Copyright 2019 Xi'an Jiaotong University

  Licensed under the Apache License, Version 2.0 (the "License");
  you may not use this file except in compliance with the License.
  You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

  Unless required by applicable law or agreed to in writing, software
  distributed under the License is distributed on an "AS IS" BASIS,
  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
  See the License for the specific language governing permissions and
  limitations under the License.
*******************************************************************************/
module LutZ3
(
	input  logic [7:0]  index,
	output logic [23:0] lut_value
);

always_comb begin
    case (index)
		8'b00000000:	lut_value = 25'b0001011001011101011001000;
		8'b00000001:	lut_value = 25'b0001011000011011011101010;
		8'b00000010:	lut_value = 25'b0001010111011010110001110;
		8'b00000011:	lut_value = 25'b0001010110011011010100101;
		8'b00000100:	lut_value = 25'b0001010101011101000011011;
		8'b00000101:	lut_value = 25'b0001010100011111111100110;
		8'b00000110:	lut_value = 25'b0001010011100011111110011;
		8'b00000111:	lut_value = 25'b0001010010101001000110001;
		8'b00001000:	lut_value = 25'b0001010001101111010010101;
		8'b00001001:	lut_value = 25'b0001010000110110100010001;
		8'b00001010:	lut_value = 25'b0001001111111110110010111;
		8'b00001011:	lut_value = 25'b0001001111001000000010111;
		8'b00001100:	lut_value = 25'b0001001110010010010001010;
		8'b00001101:	lut_value = 25'b0001001101011101011100000;
		8'b00001110:	lut_value = 25'b0001001100101001100001110;
		8'b00001111:	lut_value = 25'b0001001011110110100001010;
		8'b00010000:	lut_value = 25'b0001001011000100011000101;
		8'b00010001:	lut_value = 25'b0001001010010011000110111;
		8'b00010010:	lut_value = 25'b0001001001100010101010111;
		8'b00010011:	lut_value = 25'b0001001000110011000011001;
		8'b00010100:	lut_value = 25'b0001001000000100001110010;
		8'b00010101:	lut_value = 25'b0001000111010110001011011;
		8'b00010110:	lut_value = 25'b0001000110101000111001010;
		8'b00010111:	lut_value = 25'b0001000101111100010110100;
		8'b00011000:	lut_value = 25'b0001000101010000100010100;
		8'b00011001:	lut_value = 25'b0001000100100101011100000;
		8'b00011010:	lut_value = 25'b0001000011111011000001101;
		8'b00011011:	lut_value = 25'b0001000011010001010010110;
		8'b00011100:	lut_value = 25'b0001000010101000001110011;
		8'b00011101:	lut_value = 25'b0001000001111111110011110;
		8'b00011110:	lut_value = 25'b0001000001011000000001100;
		8'b00011111:	lut_value = 25'b0001000000110000110111000;
		8'b00100000:	lut_value = 25'b0001000000001010010011011;
		8'b00100001:	lut_value = 25'b0000111111100100010101110;
		8'b00100010:	lut_value = 25'b0000111110111110111101011;
		8'b00100011:	lut_value = 25'b0000111110011010001001011;
		8'b00100100:	lut_value = 25'b0000111101110101111001000;
		8'b00100101:	lut_value = 25'b0000111101010010001011101;
		8'b00100110:	lut_value = 25'b0000111100101111000000011;
		8'b00100111:	lut_value = 25'b0000111100001100010110011;
		8'b00101000:	lut_value = 25'b0000111011101010001101010;
		8'b00101001:	lut_value = 25'b0000111011001000100100011;
		8'b00101010:	lut_value = 25'b0000111010100111011010110;
		8'b00101011:	lut_value = 25'b0000111010000110110000000;
		8'b00101100:	lut_value = 25'b0000111001100110100011100;
		8'b00101101:	lut_value = 25'b0000111001000110110100100;
		8'b00101110:	lut_value = 25'b0000111000100111100010010;
		8'b00101111:	lut_value = 25'b0000111000001000101100101;
		8'b00110000:	lut_value = 25'b0000110111101010010010110;
		8'b00110001:	lut_value = 25'b0000110111001100010100010;
		8'b00110010:	lut_value = 25'b0000110110101110110000100;
		8'b00110011:	lut_value = 25'b0000110110010001100110111;
		8'b00110100:	lut_value = 25'b0000110101110100110111001;
		8'b00110101:	lut_value = 25'b0000110101011000100000101;
		8'b00110110:	lut_value = 25'b0000110100111100100010110;
		8'b00110111:	lut_value = 25'b0000110100100000111101010;
		8'b00111000:	lut_value = 25'b0000110100000101101111101;
		8'b00111001:	lut_value = 25'b0000110011101010111001010;
		8'b00111010:	lut_value = 25'b0000110011010000011001111;
		8'b00111011:	lut_value = 25'b0000110010110110010001000;
		8'b00111100:	lut_value = 25'b0000110010011100011110010;
		8'b00111101:	lut_value = 25'b0000110010000011000001001;
		8'b00111110:	lut_value = 25'b0000110001101001111001011;
		8'b00111111:	lut_value = 25'b0000110001010001000110011;
		8'b01000000:	lut_value = 25'b0000110000111000101000001;
		8'b01000001:	lut_value = 25'b0000110000100000011110000;
		8'b01000010:	lut_value = 25'b0000110000001000100111100;
		8'b01000011:	lut_value = 25'b0000101111110001000100100;
		8'b01000100:	lut_value = 25'b0000101111011001110100101;
		8'b01000101:	lut_value = 25'b0000101111000010110111101;
		8'b01000110:	lut_value = 25'b0000101110101100001101000;
		8'b01000111:	lut_value = 25'b0000101110010101110100011;
		8'b01001000:	lut_value = 25'b0000101101111111101101101;
		8'b01001001:	lut_value = 25'b0000101101101001111000011;
		8'b01001010:	lut_value = 25'b0000101101010100010100011;
		8'b01001011:	lut_value = 25'b0000101100111111000001001;
		8'b01001100:	lut_value = 25'b0000101100101001111110101;
		8'b01001101:	lut_value = 25'b0000101100010101001100011;
		8'b01001110:	lut_value = 25'b0000101100000000101010000;
		8'b01001111:	lut_value = 25'b0000101011101100010111101;
		8'b01010000:	lut_value = 25'b0000101011011000010100110;
		8'b01010001:	lut_value = 25'b0000101011000100100001001;
		8'b01010010:	lut_value = 25'b0000101010110000111100100;
		8'b01010011:	lut_value = 25'b0000101010011101100110101;
		8'b01010100:	lut_value = 25'b0000101010001010011111010;
		8'b01010101:	lut_value = 25'b0000101001110111100110000;
		8'b01010110:	lut_value = 25'b0000101001100100111010111;
		8'b01010111:	lut_value = 25'b0000101001010010011101101;
		8'b01011000:	lut_value = 25'b0000101001000000001110001;
		8'b01011001:	lut_value = 25'b0000101000101110001011110;
		8'b01011010:	lut_value = 25'b0000101000011100010110101;
		8'b01011011:	lut_value = 25'b0000101000001010101110011;
		8'b01011100:	lut_value = 25'b0000100111111001010011000;
		8'b01011101:	lut_value = 25'b0000100111101000000100001;
		8'b01011110:	lut_value = 25'b0000100111010111000001100;
		8'b01011111:	lut_value = 25'b0000100111000110001011001;
		8'b01100000:	lut_value = 25'b0000100110110101100000110;
		8'b01100001:	lut_value = 25'b0000100110100101000010001;
		8'b01100010:	lut_value = 25'b0000100110010100101111001;
		8'b01100011:	lut_value = 25'b0000100110000100100111100;
		8'b01100100:	lut_value = 25'b0000100101110100101011001;
		8'b01100101:	lut_value = 25'b0000100101100100111001111;
		8'b01100110:	lut_value = 25'b0000100101010101010011100;
		8'b01100111:	lut_value = 25'b0000100101000101110111111;
		8'b01101000:	lut_value = 25'b0000100100110110100111000;
		8'b01101001:	lut_value = 25'b0000100100100111100000011;
		8'b01101010:	lut_value = 25'b0000100100011000100100000;
		8'b01101011:	lut_value = 25'b0000100100001001110001110;
		8'b01101100:	lut_value = 25'b0000100011111011001001100;
		8'b01101101:	lut_value = 25'b0000100011101100101011000;
		8'b01101110:	lut_value = 25'b0000100011011110010110011;
		8'b01101111:	lut_value = 25'b0000100011010000001011001;
		8'b01110000:	lut_value = 25'b0000100011000010001001011;
		8'b01110001:	lut_value = 25'b0000100010110100010000111;
		8'b01110010:	lut_value = 25'b0000100010100110100001011;
		8'b01110011:	lut_value = 25'b0000100010011000111011001;
		8'b01110100:	lut_value = 25'b0000100010001011011101100;
		8'b01110101:	lut_value = 25'b0000100001111110001000110;
		8'b01110110:	lut_value = 25'b0000100001110000111100101;
		8'b01110111:	lut_value = 25'b0000100001100011111000111;
		8'b01111000:	lut_value = 25'b0000100001010110111101101;
		8'b01111001:	lut_value = 25'b0000100001001010001010101;
		8'b01111010:	lut_value = 25'b0000100000111101011111111;
		8'b01111011:	lut_value = 25'b0000100000110000111101000;
		8'b01111100:	lut_value = 25'b0000100000100100100010001;
		8'b01111101:	lut_value = 25'b0000100000011000001111001;
		8'b01111110:	lut_value = 25'b0000100000001100000011110;
		8'b01111111:	lut_value = 25'b0000100000000000000000000;
		8'b10000000:	lut_value = 25'b0011111010000111010111101;
		8'b10000001:	lut_value = 25'b0011111010000111010111101;
		8'b10000010:	lut_value = 25'b0011110100011100111100101;
		8'b10000011:	lut_value = 25'b0011110100011100111100101;
		8'b10000100:	lut_value = 25'b0011101110111111111111101;
		8'b10000101:	lut_value = 25'b0011101110111111111111101;
		8'b10000110:	lut_value = 25'b0011101001101111110100110;
		8'b10000111:	lut_value = 25'b0011101001101111110100110;
		8'b10001000:	lut_value = 25'b0011100100101011110010110;
		8'b10001001:	lut_value = 25'b0011100100101011110010110;
		8'b10001010:	lut_value = 25'b0011011111110011010010011;
		8'b10001011:	lut_value = 25'b0011011111110011010010011;
		8'b10001100:	lut_value = 25'b0011011011000101110000010;
		8'b10001101:	lut_value = 25'b0011011011000101110000010;
		8'b10001110:	lut_value = 25'b0011010110100010101001110;
		8'b10001111:	lut_value = 25'b0011010110100010101001110;
		8'b10010000:	lut_value = 25'b0011010010001001011110110;
		8'b10010001:	lut_value = 25'b0011010010001001011110110;
		8'b10010010:	lut_value = 25'b0011001101111001110010000;
		8'b10010011:	lut_value = 25'b0011001101111001110010000;
		8'b10010100:	lut_value = 25'b0011001001110011000110101;
		8'b10010101:	lut_value = 25'b0011001001110011000110101;
		8'b10010110:	lut_value = 25'b0011000101110101000010110;
		8'b10010111:	lut_value = 25'b0011000101110101000010110;
		8'b10011000:	lut_value = 25'b0011000001111111001100111;
		8'b10011001:	lut_value = 25'b0011000001111111001100111;
		8'b10011010:	lut_value = 25'b0010111110010001001101111;
		8'b10011011:	lut_value = 25'b0010111110010001001101111;
		8'b10011100:	lut_value = 25'b0010111010101010101111000;
		8'b10011101:	lut_value = 25'b0010111010101010101111000;
		8'b10011110:	lut_value = 25'b0010110111001011011100001;
		8'b10011111:	lut_value = 25'b0010110111001011011100001;
		8'b10100000:	lut_value = 25'b0010110011110011000000010;
		8'b10100001:	lut_value = 25'b0010110011110011000000010;
		8'b10100010:	lut_value = 25'b0010110000100001001001110;
		8'b10100011:	lut_value = 25'b0010110000100001001001110;
		8'b10100100:	lut_value = 25'b0010101101010101100110110;
		8'b10100101:	lut_value = 25'b0010101101010101100110110;
		8'b10100110:	lut_value = 25'b0010101010010000000110010;
		8'b10100111:	lut_value = 25'b0010101010010000000110010;
		8'b10101000:	lut_value = 25'b0010100111010000011000001;
		8'b10101001:	lut_value = 25'b0010100111010000011000001;
		8'b10101010:	lut_value = 25'b0010100100010110001110000;
		8'b10101011:	lut_value = 25'b0010100100010110001110000;
		8'b10101100:	lut_value = 25'b0010100001100001011001010;
		8'b10101101:	lut_value = 25'b0010100001100001011001010;
		8'b10101110:	lut_value = 25'b0010011110110001101100000;
		8'b10101111:	lut_value = 25'b0010011110110001101100000;
		8'b10110000:	lut_value = 25'b0010011100000110111001110;
		8'b10110001:	lut_value = 25'b0010011100000110111001110;
		8'b10110010:	lut_value = 25'b0010011001100000110110100;
		8'b10110011:	lut_value = 25'b0010011001100000110110100;
		8'b10110100:	lut_value = 25'b0010010110111111010110101;
		8'b10110101:	lut_value = 25'b0010010110111111010110101;
		8'b10110110:	lut_value = 25'b0010010100100010001110011;
		8'b10110111:	lut_value = 25'b0010010100100010001110011;
		8'b10111000:	lut_value = 25'b0010010010001001010011111;
		8'b10111001:	lut_value = 25'b0010010010001001010011111;
		8'b10111010:	lut_value = 25'b0010001111110100011101000;
		8'b10111011:	lut_value = 25'b0010001111110100011101000;
		8'b10111100:	lut_value = 25'b0010001101100011100000010;
		8'b10111101:	lut_value = 25'b0010001101100011100000010;
		8'b10111110:	lut_value = 25'b0010001011010110010100011;
		8'b10111111:	lut_value = 25'b0010001011010110010100011;
		8'b11000000:	lut_value = 25'b0010001001001100110000101;
		8'b11000001:	lut_value = 25'b0010001001001100110000101;
		8'b11000010:	lut_value = 25'b0010000111000110101101001;
		8'b11000011:	lut_value = 25'b0010000111000110101101001;
		8'b11000100:	lut_value = 25'b0010000101000100000001111;
		8'b11000101:	lut_value = 25'b0010000101000100000001111;
		8'b11000110:	lut_value = 25'b0010000011000100100110110;
		8'b11000111:	lut_value = 25'b0010000011000100100110110;
		8'b11001000:	lut_value = 25'b0010000001001000010101011;
		8'b11001001:	lut_value = 25'b0010000001001000010101011;
		8'b11001010:	lut_value = 25'b0001111111001111000110001;
		8'b11001011:	lut_value = 25'b0001111111001111000110001;
		8'b11001100:	lut_value = 25'b0001111101011000110011000;
		8'b11001101:	lut_value = 25'b0001111101011000110011000;
		8'b11001110:	lut_value = 25'b0001111011100101010101001;
		8'b11001111:	lut_value = 25'b0001111011100101010101001;
		8'b11010000:	lut_value = 25'b0001111001110100100111010;
		8'b11010001:	lut_value = 25'b0001111001110100100111010;
		8'b11010010:	lut_value = 25'b0001111000000110100010101;
		8'b11010011:	lut_value = 25'b0001111000000110100010101;
		8'b11010100:	lut_value = 25'b0001110110011011000010100;
		8'b11010101:	lut_value = 25'b0001110110011011000010100;
		8'b11010110:	lut_value = 25'b0001110100110010000001001;
		8'b11010111:	lut_value = 25'b0001110100110010000001001;
		8'b11011000:	lut_value = 25'b0001110011001011011001111;
		8'b11011001:	lut_value = 25'b0001110011001011011001111;
		8'b11011010:	lut_value = 25'b0001110001100111000111001;
		8'b11011011:	lut_value = 25'b0001110001100111000111001;
		8'b11011100:	lut_value = 25'b0001110000000101000100111;
		8'b11011101:	lut_value = 25'b0001110000000101000100111;
		8'b11011110:	lut_value = 25'b0001101110100101001110010;
		8'b11011111:	lut_value = 25'b0001101110100101001110010;
		8'b11100000:	lut_value = 25'b0001101101000111011111000;
		8'b11100001:	lut_value = 25'b0001101101000111011111000;
		8'b11100010:	lut_value = 25'b0001101011101011110011000;
		8'b11100011:	lut_value = 25'b0001101011101011110011000;
		8'b11100100:	lut_value = 25'b0001101010010010000110011;
		8'b11100101:	lut_value = 25'b0001101010010010000110011;
		8'b11100110:	lut_value = 25'b0001101000111010010101001;
		8'b11100111:	lut_value = 25'b0001101000111010010101001;
		8'b11101000:	lut_value = 25'b0001100111100100011011111;
		8'b11101001:	lut_value = 25'b0001100111100100011011111;
		8'b11101010:	lut_value = 25'b0001100110010000010110100;
		8'b11101011:	lut_value = 25'b0001100110010000010110100;
		8'b11101100:	lut_value = 25'b0001100100111110000010011;
		8'b11101101:	lut_value = 25'b0001100100111110000010011;
		8'b11101110:	lut_value = 25'b0001100011101101011011100;
		8'b11101111:	lut_value = 25'b0001100011101101011011100;
		8'b11110000:	lut_value = 25'b0001100010011110011111000;
		8'b11110001:	lut_value = 25'b0001100010011110011111000;
		8'b11110010:	lut_value = 25'b0001100001010001001001111;
		8'b11110011:	lut_value = 25'b0001100001010001001001111;
		8'b11110100:	lut_value = 25'b0001100000000101011001000;
		8'b11110101:	lut_value = 25'b0001100000000101011001000;
		8'b11110110:	lut_value = 25'b0001011110111011001001111;
		8'b11110111:	lut_value = 25'b0001011110111011001001111;
		8'b11111000:	lut_value = 25'b0001011101110010011001011;
		8'b11111001:	lut_value = 25'b0001011101110010011001011;
		8'b11111010:	lut_value = 25'b0001011100101011000101010;
		8'b11111011:	lut_value = 25'b0001011100101011000101010;
		8'b11111100:	lut_value = 25'b0001011011100101001010111;
		8'b11111101:	lut_value = 25'b0001011011100101001010111;
		8'b11111110:	lut_value = 25'b0001011010100000100111011;
		8'b11111111:	lut_value = 25'b0001011010100000100111011;
	endcase
end

endmodule
